module TB_v5c_sm();
  initial begin
    $display("PASSED");
    $finish;
  end
endmodule

